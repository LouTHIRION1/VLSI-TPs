library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Reg is
  port
  (
    ---- Write interface
    -- Write Port 1 prioritaire (EXEC stage)
    wdata1 : in std_logic_vector(31 downto 0);
    wadr1  : in std_logic_vector(3 downto 0); -- Register address (0 - 16)
    wen1   : in std_logic;                    -- Enable port

    -- Write Port 2 non prioritaire (MEM stage)
    wdata2 : in std_logic_vector(31 downto 0);
    wadr2  : in std_logic_vector(3 downto 0); -- Register address (0 - 16)
    wen2   : in std_logic;                    -- Enable port

    -- Write CSPR (Current Program Status Register) Port
    wneg    : in std_logic; -- Write N flag
    wzero   : in std_logic; -- Write Z flag
    wcry    : in std_logic; -- Write C flag
    wovr    : in std_logic; -- Write V flag
    cpsr_wb : in std_logic; -- CPSR register writeback enable

    ---- Read interface
    -- Read Port 1 32 bits (Rd)
    reg_rd1 : out std_logic_vector(31 downto 0); -- Register 1
    radr1   : in std_logic_vector(3 downto 0);   -- Register 1 address (0 - 16)
    reg_v1  : out std_logic;                     -- Register 1 validity bit

    -- Read Port 2 32 bits (Rs)
    reg_rd2 : out std_logic_vector(31 downto 0); -- Register 2
    radr2   : in std_logic_vector(3 downto 0);   -- Register 2 address (0 - 16)
    reg_v2  : out std_logic;                     -- Register 2 validity bit

    -- Read Port 3 32 bits (Rt)
    reg_rd3 : out std_logic_vector(31 downto 0); -- Register 3
    radr3   : in std_logic_vector(3 downto 0);   -- Register 3 address (0 - 16)
    reg_v3  : out std_logic;                     -- Register 3 validity bit

    ---- CPSR
    -- Read CPSR (Current Program Status Register) Port
    reg_neg  : out std_logic; -- Read N flag
    reg_zero : out std_logic; -- Read Z flag
    reg_cry  : out std_logic; -- Read C flag
    reg_cznv : out std_logic; -- CZN flag validity (for logic instructions)
    reg_ovr  : out std_logic; -- Read V flag
    reg_vv   : out std_logic; -- V flag validity(for arithmetic instructions)

    ---- Invalidation
    -- Invalidate Port 1
    inval_adr1 : in std_logic_vector(3 downto 0); -- Invalidate address Register 1 (0 - 16)
    inval1     : in std_logic;                    -- Invalidate Register 1
    -- Invalidate Port 2
    inval_adr2 : in std_logic_vector(3 downto 0); -- Invalidate address Register 2 (0 - 16)
    inval2     : in std_logic;                    -- Invalidate Register 2
    -- Invalidate Flags
    inval_czn : in std_logic; -- Invalidate C Z N flags (Logic instructions)
    inval_ovr : in std_logic; -- Invalidate V flag (Arithmetic instructions)

    ---- Program Counter (PC)
    reg_pc  : out std_logic_vector(31 downto 0); -- Program Counter register
    reg_pcv : out std_logic;                     -- Program Counter validity
    inc_pc  : in std_logic;                      -- Increment PC +4

    -- global interface
    clk     : in std_logic; -- Clock
    reset_n : in std_logic; -- Reset (active low)
    vdd     : in bit;
    vss     : in bit);
end Reg;

architecture behavioral_reg of Reg is
  -- Registers 1 - 12
  signal registre0  : std_logic_vector(31 downto 0);
  signal registre1  : std_logic_vector(31 downto 0);
  signal registre2  : std_logic_vector(31 downto 0);
  signal registre3  : std_logic_vector(31 downto 0);
  signal registre4  : std_logic_vector(31 downto 0);
  signal registre5  : std_logic_vector(31 downto 0);
  signal registre6  : std_logic_vector(31 downto 0);
  signal registre7  : std_logic_vector(31 downto 0);
  signal registre8  : std_logic_vector(31 downto 0);
  signal registre9  : std_logic_vector(31 downto 0);
  signal registre10 : std_logic_vector(31 downto 0);
  signal registre11 : std_logic_vector(31 downto 0);
  signal registre12 : std_logic_vector(31 downto 0);
  -- Register SP
  signal registre13 : std_logic_vector(31 downto 0);
  -- Register LR
  signal registre14 : std_logic_vector(31 downto 0);
  -- Register PC
  signal registre15 : std_logic_vector(31 downto 0);

  signal CPSR : std_logic_vector(3 downto 0);

begin
  process (clk)
  begin
    -- Synchronous
    if rising_edge(clk) then
      if (reset_n = '0') then
        -- Invalidate Register ports
        reg_v1 <= '1';
        reg_v2 <= '1';
        reg_v3 <= '1';
        -- Reset CPSR
        reg_cry  <= '0'; -- C fag
        reg_zero <= '0'; -- Z flag
        reg_neg  <= '0'; -- N flag
        reg_ovr  <= '0'; -- V flag
        reg_cznv <= '0'; -- CZN Validity bit (arithmetic)
        reg_vv   <= '0'; -- V Validity bit (logic)
      else
        -- Write CPSR register when writeback is enabled
        if (cpsr_wb = '1') then
          -- N flag
          reg_neg <= wneg when (reg_cznv_s = '1') else
            reg_neg;
          -- Z flag
          reg_zero <= wzero when (reg_cznv_s = '1') else
            reg_zero;
          -- C flag
          reg_cry <= wcry when (reg_cznv_s = '1') else
            reg_cry;
          -- V flag
          reg_ovr <= wovr when (reg_vv_s = '1') else
            reg_ovr;

        end if;
      end if;
    end if;
  end process;
end behavioral_reg;
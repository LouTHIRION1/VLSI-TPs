* description d'un inverseur CMOS

.lib typical
.include ../mosn_mosp.wc
.lib "mon_inv.spi" circuit
.endl  typical

.lib circuit
.subckt mon_inv d q vdd vss bn bp param: W=2.0e-06
MP q d vdd bp TP L=0.35e-06 W=W
MN q d vss bn TN L=0.35e-06 W=1.4e-06
.ends

.endl circuit
